module alu(
    input logic clk,
    input logic rst,
    input logic dump // 用于控制波形记录
);
    // 其他逻辑...
endmodule
